library IEEE;
use IEEE.STD_LOGIC_1164.all;

package Common_Types_Pck is

	type buscar is array (0 to 10) of STD_LOGIC_VECTOR(20 downto 1);

end Common_Types_Pck;